--Alan Decowski
--CPE 487
--2021F
--font.vhd
--ACCEPTS: char
--Char: An integer that references a bitmap within character set.

--RETURNS: bits
--bits: a 64-bit word containing the bitmap of the requested character code.

library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.std_logic_arith.ALL;


entity font is
 Port ( 
 char : IN integer;
 bits : OUT std_logic_vector(63 DOWNTO 0)
 );
end font;

architecture Behavioral of font is
begin
		bits <= "0000000000000000000000000000000000000000000000000000000000000000" WHEN char = 0 ELSE -- 
				"0000000000011000001001000100001001000010011111100100001001000010" WHEN char = 1 ELSE --A
				"0000000001111100010000100100001001111100010000100100001001111100" WHEN char = 2 ELSE --B
				"0000000000111110010000000100000001000000010000000100000000111110" WHEN char = 3 ELSE --C
				"0000000001111000010001000100001001000010010000100100010001111000" WHEN char = 4 ELSE --D
				"0000000001111110010000000100000001111100010000000100000001111110" WHEN char = 5 ELSE --E
				"0000000001111110010000000100000001111100010000000100000001000000" WHEN char = 6 ELSE --F
				"0000000001111110010000000100000001011110010000100100001001111110" WHEN char = 7 ELSE --G
				"0000000001000010010000100100001001111110010000100100001001000010" WHEN char = 8 ELSE --H
				"0000000011111110000100000001000000010000000100000001000011111110" WHEN char = 9 ELSE --I
				"0000000011111110000100000001000000010000000100000001000011100000" WHEN char = 10 ELSE --J
				"0000000001000010010001000101100001100000010110000100010001000010" WHEN char = 11 ELSE --K
				"0000000001000000010000000100000001000000010000000100000001111100" WHEN char = 12 ELSE --L
				"0000000011000110101010101001001010010010100100101001001010010010" WHEN char = 13 ELSE --M
				"0000000001100010010100100101001001001010010010100100011001000110" WHEN char = 14 ELSE --N
				"0000000000111000010001001000001010000010100000100100010000111000" WHEN char = 15 ELSE --O
				"0000000001111000010001000100010001111000010000000100000001000000" WHEN char = 16 ELSE --P
				"0000000000111000010001001000001010000010100010100100010000111010" WHEN char = 17 ELSE --Q
				"0000000001111100010000100100001001111100010000100100001001000010" WHEN char = 18 ELSE --R
				"0000000000111110010000000100000000111100000000100000001001111100" WHEN char = 19 ELSE --S
				"0000000011111110000100000001000000010000000100000001000000010000" WHEN char = 20 ELSE --T
				"0000000001000010010000100100001001000010010000100100001000111100" WHEN char = 21 ELSE --U
				"0000000001000010010000100100001001000010010000100010010000011000" WHEN char = 22 ELSE --V
				"0000000010010010100100101001001010010010100100101010101011000110" WHEN char = 23 ELSE --W
				"0000000010000010010001000010100000010000001010000100010010000010" WHEN char = 24 ELSE --X
				"0000000001000100010001000010100000101000000100000001000000010000" WHEN char = 25 ELSE --Y
				"0000000011111100000011000001000000100000010000001000000011111100" WHEN char = 26 ELSE --Z
				"0000000000010000001100000101000000010000000100000001000001111100" WHEN char = 27 ELSE --1
				"0000000000111000010001000000010000001000000100000010000001111100" WHEN char = 28 ELSE --2
				"0000000001111000000001000000010001111000000001000000010001111000" WHEN char = 29 ELSE --3
				"0000000001000100010001000100010001111100000001000000010000000100" WHEN char = 30 ELSE --4
				"0000000001111100010000000100000001111100000001000100010000111000" WHEN char = 31 ELSE --5
				"0000000000111110010000000100000001111100010000100100001000111100" WHEN char = 32 ELSE --6
				"0000000001111110000000100000010000001000000100000010000001000000" WHEN char = 33 ELSE --7
				"0000000000111100010000100100001000111100010000100100001000111100" WHEN char = 34 ELSE --8
				"0000000000111000010001000100010000111100000001000000010001111000" WHEN char = 35 ELSE --9
				"0000000001111100100001101000101010010010101000101100001001111100" WHEN char = 36 ELSE --0
				"0000000000011000000110000000000000000000000110000001100000000000" WHEN char = 37 ELSE --:
				"0000000000000000000000000000000000000000000000000000000000000000";

end Behavioral;
